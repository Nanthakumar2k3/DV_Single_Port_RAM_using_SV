`include "memory.sv"
`include "common.sv"
`include "mem_intf.sv"
`include "mem_tx.sv"
`include "mem_gen.sv"
`include "mem_bfm.sv"
`include "mem_mon.sv"
`include "mem_cov.sv"
`include "mem_agent.sv"
`include "mem_sbd.sv"
`include "mem_env.sv"
`include "top.sv"


// typedef class mem_gen;
// typedef class mem_bfm;
// typedef class mem_mon;
// typedef class mem_cov;
// typedef class mem_sbd;
// typedef class mem_agent;
// typedef class mem_env;


// `include "mem_gen.sv"
// `include "mem_cov.sv"
// `include "mem_bfm.sv"
// `include "mem_mon.sv"
// `include "mem_env.sv"
// `include "mem_agent.sv"
// `include "mem_sbd.sv"
// `include "top.sv"








